,src_ip,,AS13335 CLOUDFLARENET,AS13414 TWITTER,AS14061 DIGITALOCEAN-ASN,AS14618 AMAZON-AES,AS14907 WIKIMEDIA,AS15169 GOOGLE,AS15525 Servicos De Comunicacoes E Multimedia S.A.,AS16509 AMAZON-02,AS16625 AKAMAI-AS,"AS1930 Fundacao para a Ciencia e a Tecnologia, I.P.",AS19551 INCAPSULA,AS20940 Akamai International B.V.,AS24768 Almouroltec Servicos De Informatica E Internet Lda,AS24940 Hetzner Online GmbH,"AS2860 Nos Comunicacoes, S.A.",AS29789 REFLECTED,AS31898 ORACLE-BMC-31898,AS32244 LIQUIDWEB,AS3243 Servicos De Comunicacoes E Multimedia S.A.,AS32934 FACEBOOK,AS35995 TWITTER,AS36459 GITHUB,AS396982 GOOGLE-CLOUD-PLATFORM,AS43515 Google Ireland Limited,AS46652 SERVERSTACK-ASN,AS54113 FASTLY,AS54115 FACEBOOK-CORP,AS6167 CELLCO-PART,AS62540 DRAKE-AS,AS62785 AMAZON-FC,AS63179 TWITTER,AS63194 CRASH,AS63949 Akamai Connected Cloud,AS7018 ATT-INTERNET4,AS7224 AMAZON-AS,AS8068 MICROSOFT-CORP-MSN-AS-BLOCK,AS8069 MICROSOFT-CORP-MSN-AS-BLOCK,AS8070 MICROSOFT-CORP-MSN-AS-BLOCK,AS8075 MICROSOFT-CORP-MSN-AS-BLOCK,AS8657 Servicos De Comunicacoes E Multimedia S.A.,AS8987 Amazon Data Services Ireland Ltd,"AS9186 Infocomunicacoes, S.A."
44,192.168.107.140,4336,343,340,65,26,253,1713,406,56,12,114,1,2,1,248,1071,128,126,34,510,1447,4,0,31,14,205,109,0,0,0,0,0,0,110,0,3,393,0,3,452,45,0,65
150,192.168.107.51,4176,202,262,12,6,208,1631,301,107,16,21,6,23,9,192,943,117,67,44,506,1283,2,0,20,5,254,101,4,0,4,6,12,14,165,0,0,425,0,91,433,22,3,46
42,192.168.107.139,4007,346,392,34,10,286,1780,286,68,7,77,15,4,58,285,848,105,130,21,378,1191,0,0,16,0,180,109,0,0,0,0,0,0,152,2,0,419,0,17,399,43,0,93
169,192.168.107.70,3610,181,251,28,12,240,1648,301,65,6,38,22,4,1,226,762,65,131,8,475,1258,0,0,16,0,195,69,0,0,0,0,0,0,85,2,0,361,0,34,392,50,0,86
41,192.168.107.138,3606,342,308,49,4,166,1460,195,84,7,48,12,0,6,144,818,64,66,61,429,904,0,0,18,0,155,113,0,0,0,0,0,0,133,8,0,326,0,32,400,35,0,36
145,192.168.107.46,3559,256,301,38,42,278,1572,220,66,3,70,9,0,11,288,856,114,63,11,496,1032,2,2,38,0,271,50,0,0,0,3,0,0,187,0,5,337,0,9,353,29,0,102
62,192.168.107.157,3497,168,293,21,30,190,1346,179,46,4,88,6,0,0,183,619,64,105,29,509,1275,0,0,16,0,128,101,0,0,8,0,0,0,139,0,17,395,0,56,392,14,0,27
119,192.168.107.21,3482,337,379,34,10,279,1392,221,45,10,82,26,13,3,136,780,31,50,14,482,1332,0,0,6,0,288,104,0,0,0,0,3,0,150,2,0,313,0,47,274,10,0,143
91,192.168.107.184,3467,310,287,66,10,270,1592,183,60,34,98,5,0,0,222,644,90,38,47,429,899,0,0,15,0,137,25,0,0,0,0,20,0,92,0,0,281,0,22,316,35,0,24
26,192.168.107.124,3448,199,247,11,0,265,1428,243,42,0,71,0,3,23,152,920,71,59,23,373,988,0,4,6,18,135,55,0,0,0,0,8,0,116,0,0,367,0,97,330,41,1,38
179,192.168.107.80,3446,250,344,43,5,218,1431,281,115,4,51,14,2,5,216,930,95,75,10,467,1046,2,0,22,0,202,118,1,0,0,0,1,2,169,6,0,370,0,6,273,34,0,15
146,192.168.107.47,3440,252,341,32,0,155,1511,172,52,20,64,12,6,18,116,862,39,82,8,370,1142,7,0,29,0,179,76,1,0,0,3,0,0,72,0,0,292,0,16,333,44,0,41
89,192.168.107.182,3432,269,285,31,11,193,1397,231,38,0,47,3,0,11,146,718,80,69,18,415,1088,5,1,27,0,166,104,0,0,0,6,0,0,103,0,0,393,0,24,351,13,2,49
104,192.168.107.196,3406,321,297,40,0,171,1496,155,35,5,35,1,7,0,202,726,72,92,41,345,1011,12,8,31,1,193,85,0,0,0,0,0,0,103,0,3,242,0,9,294,14,0,26
7,192.168.107.107,3369,248,239,23,23,170,1463,252,98,4,54,29,12,0,208,737,70,92,15,443,993,1,3,16,0,123,115,0,0,4,0,0,0,91,8,13,355,2,4,402,13,0,30
88,192.168.107.181,3326,357,231,51,1,174,1349,194,55,24,65,21,10,2,230,874,92,109,5,446,1096,0,0,49,0,192,118,0,0,0,1,0,0,123,0,5,342,0,1,281,66,0,56
152,192.168.107.53,3186,283,260,25,21,298,1335,195,40,0,80,7,8,0,174,684,48,96,33,405,1040,0,0,14,0,153,139,0,1,0,0,12,4,179,1,0,358,0,19,270,17,0,76
117,192.168.107.208,3164,250,217,34,11,201,1443,176,65,23,46,10,16,8,170,737,99,142,78,408,964,0,0,8,0,125,31,0,0,0,6,0,0,89,0,6,287,0,35,276,52,0,77
50,192.168.107.146,3090,214,291,21,2,209,1386,144,31,8,19,0,9,0,222,714,44,65,7,313,898,0,4,39,0,172,102,0,0,0,5,0,7,156,0,0,350,0,33,288,31,0,33
138,192.168.107.39,3076,261,294,16,2,176,1342,214,85,5,44,5,8,0,190,539,115,111,19,444,949,5,0,42,0,192,54,0,0,0,3,0,0,207,16,0,281,0,41,424,48,0,25
184,192.168.107.85,2969,308,299,27,13,169,1471,174,34,12,59,4,11,16,172,816,87,82,37,471,881,4,0,24,0,215,88,0,0,0,0,3,0,102,0,3,356,0,7,362,8,0,119
137,192.168.107.38,2943,356,279,17,2,178,1342,180,71,23,51,4,0,0,111,676,72,122,17,324,918,0,0,27,10,136,61,0,0,0,2,1,0,61,0,0,237,0,14,266,18,0,54
191,192.168.107.92,2887,208,303,13,21,155,1172,231,45,8,58,6,25,0,218,504,150,85,13,252,888,0,0,8,0,211,73,0,0,0,12,0,0,105,7,0,239,0,35,341,1,0,33
101,192.168.107.193,2816,147,280,45,1,122,1018,176,62,9,52,12,7,0,147,608,60,75,8,451,922,1,0,9,0,207,61,0,0,0,0,2,0,95,12,0,285,0,37,285,6,0,58
190,192.168.107.91,2757,239,281,73,15,128,1161,229,49,7,45,1,23,1,189,449,60,84,30,318,895,0,0,35,0,152,73,0,0,1,3,0,0,122,4,0,312,0,14,275,49,0,25
124,192.168.107.25,2756,204,178,3,1,199,1147,151,44,0,90,9,0,9,116,725,88,73,16,425,762,3,0,0,0,117,62,7,0,0,0,0,0,87,0,3,173,0,17,263,13,2,30
114,192.168.107.205,2745,168,259,17,29,170,1026,256,81,0,35,5,0,14,111,870,50,84,18,348,837,0,1,19,0,59,82,0,0,0,0,0,0,62,0,14,259,0,5,187,34,0,44
167,192.168.107.68,2738,249,218,12,19,165,1074,189,81,1,46,3,5,0,174,748,103,130,5,291,819,0,9,10,0,112,68,0,0,3,0,0,0,105,0,0,333,0,15,341,25,0,54
72,192.168.107.167,2723,272,242,19,6,150,1256,172,54,1,65,2,9,1,86,536,52,84,51,430,900,0,0,34,0,183,127,0,0,0,0,15,0,106,0,0,246,0,27,296,20,0,54
131,192.168.107.32,2649,146,220,20,8,118,853,200,64,4,47,40,0,4,93,574,19,70,13,326,840,0,0,24,0,166,65,0,0,0,0,0,0,77,7,0,233,0,1,281,24,0,44
143,192.168.107.44,2647,239,215,35,13,152,1352,225,30,13,28,13,0,2,173,579,72,50,6,341,827,0,0,9,0,208,57,0,0,0,0,0,0,119,0,0,297,0,27,291,10,0,50
197,192.168.107.98,2624,234,247,17,13,200,1251,202,38,10,6,20,0,10,185,674,99,39,5,397,638,0,0,14,3,167,51,0,4,0,0,7,0,58,0,4,375,0,7,338,17,0,31
4,192.168.107.104,2570,183,204,18,0,138,1104,116,68,6,50,1,3,1,130,603,73,42,14,234,926,0,0,19,0,108,68,0,0,0,7,0,0,80,0,1,223,0,15,302,5,0,36
160,192.168.107.61,2555,132,212,29,14,208,999,215,64,0,27,0,10,0,191,553,73,81,9,298,883,6,0,21,0,161,39,0,0,0,0,1,8,104,0,0,293,0,29,240,17,0,50
144,192.168.107.45,2529,293,137,4,0,107,1136,161,22,4,62,3,0,0,111,593,62,25,20,327,738,3,0,18,0,164,69,0,4,0,0,0,0,52,2,3,241,0,0,230,1,0,42
10,192.168.107.11,2521,151,229,41,13,125,979,134,98,4,22,2,0,0,142,548,36,44,18,210,837,0,0,28,0,181,39,1,0,0,13,0,0,114,0,0,235,0,6,227,4,0,75
95,192.168.107.188,2512,266,231,11,21,148,1032,152,24,0,31,10,0,12,94,559,71,53,0,310,791,14,0,19,0,150,20,7,0,1,0,3,0,65,0,0,228,0,14,388,5,0,66
111,192.168.107.202,2505,195,169,30,3,148,1274,210,59,0,59,3,0,0,129,607,70,58,45,347,882,0,0,2,0,172,80,0,0,0,0,2,0,99,11,0,261,0,11,330,37,0,91
175,192.168.107.76,2465,173,252,14,5,122,1317,212,63,1,112,1,0,9,158,538,31,50,25,278,953,1,0,15,0,205,64,0,0,0,8,2,0,63,0,0,276,0,26,267,22,0,30
18,192.168.107.117,2459,187,183,5,3,130,1034,182,61,4,36,19,0,0,82,515,49,85,0,196,685,0,0,41,0,138,35,0,0,0,0,0,0,80,0,0,187,0,38,227,28,0,26
128,192.168.107.29,2448,214,244,32,1,123,1065,160,36,1,48,10,1,0,228,767,61,35,50,309,841,0,0,64,0,120,45,0,0,0,0,0,0,78,2,0,222,0,16,273,10,0,29
174,192.168.107.75,2413,244,352,19,28,184,1015,162,65,13,67,13,1,23,125,525,44,55,9,303,779,0,0,15,0,221,45,0,0,0,0,0,0,95,0,0,220,0,20,210,13,0,17
136,192.168.107.37,2408,210,160,7,0,138,1007,166,28,0,77,0,0,0,102,571,40,65,26,261,799,2,0,8,0,90,77,0,0,3,0,2,0,48,0,4,257,0,7,334,26,0,70
70,192.168.107.164,2403,90,170,11,0,101,980,178,51,4,47,1,0,7,154,565,43,46,1,233,710,0,0,9,0,104,62,0,0,0,6,0,0,64,0,0,257,0,28,251,8,0,34
192,192.168.107.93,2373,223,244,30,0,142,991,121,28,2,45,0,0,2,114,570,27,40,8,317,640,0,0,7,0,144,65,0,0,0,0,2,0,62,0,0,167,0,19,200,8,0,24
103,192.168.107.195,2350,183,189,19,22,155,1056,158,62,0,64,0,13,0,116,496,50,73,53,342,668,9,0,22,0,111,46,2,0,0,0,0,0,162,0,0,191,0,4,180,34,0,78
30,192.168.107.128,2332,188,145,14,5,120,1150,338,109,10,28,0,4,0,108,557,56,60,15,335,683,0,0,11,3,142,62,5,0,0,1,1,0,133,0,0,257,0,31,302,24,0,33
177,192.168.107.78,2309,135,198,8,0,155,930,99,27,0,30,17,5,2,63,498,25,38,19,276,800,3,0,39,0,130,75,6,0,0,0,0,0,87,0,0,249,0,14,174,27,0,18
173,192.168.107.74,2306,138,238,62,3,233,1363,180,17,0,7,4,9,1,104,542,45,104,24,277,848,0,0,28,5,181,67,0,0,0,0,0,0,86,0,0,186,0,26,222,19,0,16
118,192.168.107.209,2305,212,182,48,7,114,1067,143,64,0,22,2,0,6,111,513,41,101,41,305,886,35,1,17,0,120,36,0,0,0,0,0,0,110,0,0,187,0,23,235,19,0,37
96,192.168.107.189,2275,153,196,11,0,188,842,206,48,2,33,4,0,5,67,517,34,50,19,291,660,0,0,14,0,119,144,0,0,0,0,0,0,49,0,2,195,0,15,215,35,0,56
140,192.168.107.41,2268,143,164,11,18,114,1070,140,37,1,90,1,0,0,113,483,51,34,22,300,772,0,0,7,0,131,65,0,0,0,13,0,0,46,0,0,210,0,6,219,16,0,35
194,192.168.107.95,2246,111,211,22,14,141,865,206,23,10,63,3,0,2,84,470,38,45,17,255,596,0,0,4,2,139,35,0,0,0,0,0,0,80,0,0,185,0,32,248,16,0,9
78,192.168.107.172,2244,84,133,5,7,135,868,148,19,2,118,0,9,0,149,548,27,65,28,232,623,0,0,9,0,114,49,0,0,9,0,0,0,94,0,0,174,0,14,154,43,0,54
141,192.168.107.42,2234,159,181,6,26,178,982,248,71,10,44,3,20,0,85,491,51,86,27,335,641,0,0,11,0,80,22,0,0,0,0,0,0,61,0,0,252,0,32,197,25,0,33
161,192.168.107.62,2210,186,177,11,8,154,927,116,46,6,31,0,2,0,219,523,65,33,54,321,703,2,0,16,0,141,84,0,0,0,0,0,0,56,0,0,225,0,31,193,13,0,114
39,192.168.107.136,2186,188,206,12,5,192,1060,188,35,6,49,0,5,0,170,485,78,45,12,194,857,0,6,11,0,108,37,3,13,30,0,0,0,80,0,0,205,0,14,144,10,0,14
29,192.168.107.127,2184,158,168,20,6,165,1150,129,10,1,59,0,0,2,127,501,54,90,17,298,664,0,0,25,3,129,117,0,0,0,0,0,0,104,0,10,235,0,10,244,16,0,22
92,192.168.107.185,2179,156,170,11,5,179,764,113,23,0,20,0,1,3,76,484,39,37,0,311,624,0,0,17,0,107,56,0,11,0,0,0,0,98,0,0,129,0,12,184,21,0,22
64,192.168.107.159,2174,153,209,3,11,130,883,75,8,5,24,5,0,7,102,455,102,63,20,244,715,0,0,9,11,156,50,0,0,0,0,0,0,63,0,0,191,0,5,222,34,0,30
43,192.168.107.14,2173,180,154,19,5,111,839,117,21,1,32,4,0,0,162,508,64,65,62,282,669,1,0,24,15,136,35,0,0,0,1,0,0,90,0,0,122,0,34,181,4,0,46
53,192.168.107.149,2155,200,221,34,15,141,866,123,49,0,31,3,0,19,142,467,48,55,26,280,675,2,0,5,0,97,62,0,0,1,0,0,0,69,0,0,263,0,22,305,42,0,19
168,192.168.107.69,2154,242,154,24,0,148,921,159,15,8,46,8,30,5,162,594,41,30,2,244,669,0,0,8,0,125,90,0,0,0,0,0,0,64,0,0,230,0,9,207,9,0,24
36,192.168.107.133,2130,173,137,12,0,152,853,100,12,3,11,4,0,11,103,488,83,51,2,267,565,0,0,10,0,115,25,0,0,0,0,0,0,117,3,11,316,0,7,229,6,0,51
139,192.168.107.40,2123,126,199,13,6,113,888,182,39,0,51,1,0,0,111,410,21,38,11,346,585,0,0,60,0,136,65,0,0,0,0,0,0,40,0,1,171,0,18,332,4,0,27
151,192.168.107.52,2097,179,137,11,12,205,857,116,35,0,66,0,0,2,111,337,35,35,17,333,525,4,0,15,0,97,35,0,0,0,0,0,0,55,0,1,265,0,4,160,4,6,40
93,192.168.107.186,2083,108,164,31,4,83,933,70,37,14,50,0,0,12,50,566,41,38,19,232,788,2,0,9,0,138,30,0,0,0,0,0,0,96,4,0,176,0,7,261,42,0,56
195,192.168.107.96,2073,184,232,21,10,144,761,151,101,10,39,0,2,0,94,489,23,25,11,283,630,0,0,5,0,104,55,0,0,0,0,4,0,116,0,0,200,0,18,165,20,0,16
107,192.168.107.199,2064,151,186,42,17,131,1050,224,16,0,81,0,0,3,124,466,60,96,23,377,626,8,0,16,0,113,61,0,0,0,7,0,0,41,0,0,314,0,17,217,42,0,44
134,192.168.107.35,2060,144,200,27,4,149,882,192,56,0,64,0,4,0,129,369,44,83,12,342,589,0,0,15,0,103,46,0,0,0,0,0,0,107,0,0,221,0,18,235,23,0,43
33,192.168.107.130,2035,120,167,21,0,149,936,120,13,0,80,13,7,0,100,432,64,42,3,243,582,3,0,0,5,142,83,0,0,0,0,13,0,68,0,0,298,0,19,165,10,0,28
1,192.168.107.101,2029,81,167,22,6,86,822,72,53,0,65,6,0,0,79,449,74,65,5,365,557,2,0,5,0,80,37,0,0,0,0,0,0,136,5,3,158,0,11,168,0,0,41
40,192.168.107.137,2019,147,132,15,5,154,818,131,29,2,48,0,3,0,73,457,30,25,16,247,542,17,0,18,0,131,75,0,0,0,0,14,0,82,0,0,193,0,10,236,38,4,47
9,192.168.107.109,1981,115,163,0,6,117,820,126,30,0,61,17,10,1,88,497,45,28,7,226,512,0,0,24,0,75,16,0,0,0,0,0,0,53,0,0,189,0,17,222,9,0,45
32,192.168.107.13,1938,141,126,13,4,132,648,69,27,0,49,0,1,4,99,274,14,26,1,125,557,0,0,12,0,132,41,0,0,0,0,0,0,58,0,3,131,0,27,112,18,0,26
147,192.168.107.48,1937,171,145,36,4,96,777,123,28,3,43,17,2,0,104,490,25,54,1,314,615,14,0,0,0,88,71,0,0,0,15,0,0,28,0,0,201,0,39,174,7,0,33
102,192.168.107.194,1934,235,191,12,3,124,980,146,10,0,57,7,0,0,102,376,30,43,25,357,577,0,0,2,0,106,53,0,2,6,0,1,0,63,0,9,210,0,31,146,3,0,45
125,192.168.107.26,1930,148,98,12,0,150,746,121,19,1,40,0,0,0,153,350,72,34,1,145,669,0,0,23,0,56,41,0,0,0,0,0,0,103,0,0,215,0,23,144,8,1,28
100,192.168.107.192,1928,210,190,27,4,140,856,98,17,1,87,7,4,17,111,318,27,59,45,276,444,0,1,8,0,76,66,0,0,0,11,5,0,54,0,0,152,0,26,186,12,0,46
130,192.168.107.31,1928,138,291,8,0,116,895,109,47,0,64,13,0,0,90,406,28,34,13,320,704,0,0,18,0,78,19,0,0,0,0,0,0,117,0,0,146,1,11,143,37,0,33
85,192.168.107.179,1912,137,156,0,31,100,755,160,27,10,29,0,0,0,58,504,49,41,0,257,644,5,0,36,0,109,12,0,0,1,0,0,0,73,1,0,221,0,21,185,5,0,49
59,192.168.107.154,1892,254,150,23,6,124,841,89,32,1,8,3,0,10,95,453,3,35,24,291,573,0,0,12,0,133,43,0,0,0,0,0,7,74,2,0,223,0,21,114,19,0,29
71,192.168.107.166,1887,68,133,37,0,92,825,89,19,7,36,46,0,0,36,462,35,45,40,141,541,1,0,3,0,142,96,0,0,0,0,0,0,57,0,0,169,0,13,199,23,0,24
183,192.168.107.84,1867,110,216,18,21,91,883,174,26,0,55,0,5,15,145,487,89,56,62,309,662,0,0,18,0,126,50,0,3,0,0,0,0,65,0,0,244,0,11,208,8,0,53
81,192.168.107.175,1833,121,199,45,10,172,998,60,52,5,28,21,8,0,150,500,47,96,27,257,584,0,0,13,0,95,16,0,0,5,0,0,0,43,0,0,205,0,2,114,17,0,32
178,192.168.107.79,1832,124,85,0,9,109,758,131,3,3,22,4,0,13,76,449,84,72,22,256,607,0,0,19,0,148,83,0,0,1,0,0,0,76,0,0,191,0,18,181,13,0,19
3,192.168.107.103,1828,203,246,18,0,90,788,145,46,5,80,8,0,18,121,322,19,44,13,231,601,0,0,25,0,114,29,0,0,0,0,2,0,88,0,0,207,0,0,192,14,0,42
157,192.168.107.58,1822,92,191,3,21,108,717,119,42,0,52,0,0,0,149,360,36,43,5,119,442,0,2,10,0,36,51,0,0,0,0,0,0,76,0,3,146,0,6,177,7,0,9
105,192.168.107.197,1822,127,118,31,0,135,798,135,45,0,70,0,0,18,85,397,57,67,11,149,676,19,0,30,0,74,53,0,0,0,0,2,0,50,0,0,217,0,11,169,2,0,35
22,192.168.107.120,1819,131,153,0,1,173,818,98,21,6,57,22,0,6,65,401,33,36,15,179,605,1,0,7,0,134,50,0,0,0,0,0,0,53,0,0,215,0,17,193,27,2,6
55,192.168.107.150,1805,191,244,25,2,148,1014,121,44,20,47,5,0,0,62,487,46,42,2,181,595,0,6,18,0,119,45,0,0,0,0,0,0,63,0,0,149,0,5,247,9,0,31
75,192.168.107.17,1788,129,153,22,0,108,771,138,58,0,38,13,6,0,127,412,23,59,8,290,422,7,0,1,7,105,72,0,0,0,0,0,0,122,0,0,143,0,7,249,23,9,20
106,192.168.107.198,1782,142,122,31,8,143,801,99,40,1,46,4,13,6,58,404,25,77,2,210,526,18,14,6,0,116,72,0,0,0,0,18,0,70,0,0,195,0,24,209,9,0,16
112,192.168.107.203,1778,119,116,0,7,133,802,148,75,2,49,5,2,8,70,331,37,75,9,242,550,0,0,1,0,74,24,0,0,0,0,0,0,74,0,0,162,0,5,195,0,0,20
35,192.168.107.132,1758,147,150,6,0,63,691,91,42,0,43,0,0,14,63,330,48,88,19,247,511,0,9,3,0,70,47,0,0,0,0,0,0,119,0,0,248,0,6,121,9,6,14
77,192.168.107.171,1754,109,209,39,2,149,947,168,26,0,31,7,1,1,113,530,57,31,1,256,589,0,0,36,0,140,25,0,0,0,0,5,0,63,0,0,130,0,16,201,12,0,31
19,192.168.107.118,1746,144,94,9,3,64,735,97,33,2,34,3,9,0,118,426,32,18,20,179,511,7,0,4,0,106,34,0,0,0,0,12,0,87,0,0,122,0,31,132,4,0,28
21,192.168.107.12,1744,129,154,5,0,130,688,91,13,7,5,0,18,0,113,407,12,56,19,164,503,0,0,11,0,136,73,0,0,0,0,0,0,37,0,0,202,0,14,110,0,0,17
155,192.168.107.56,1738,137,159,8,0,139,879,178,25,4,74,0,0,10,132,452,51,54,17,158,464,0,0,8,2,167,13,0,0,0,0,0,0,72,0,0,179,0,0,156,36,0,47
171,192.168.107.72,1735,141,182,15,15,131,955,98,37,0,53,0,0,4,108,459,41,36,12,310,509,0,0,17,0,100,43,0,0,0,0,0,0,71,0,6,191,0,11,80,0,0,35
148,192.168.107.49,1732,108,193,3,2,161,792,102,23,2,57,7,0,2,57,457,74,67,9,243,590,0,0,13,0,74,83,0,0,0,0,0,0,77,0,14,146,0,1,177,12,2,0
129,192.168.107.30,1718,137,215,0,6,129,656,117,69,0,44,3,4,7,95,489,32,43,10,325,592,0,0,13,0,171,31,0,0,0,0,0,6,76,0,0,197,0,2,103,7,0,28
159,192.168.107.60,1716,116,163,11,8,92,812,72,65,0,81,0,5,0,62,363,59,14,29,141,614,0,0,8,0,126,30,0,0,3,0,0,2,41,0,0,151,0,6,146,6,0,11
164,192.168.107.65,1711,119,197,24,0,87,839,115,17,0,42,2,0,0,110,365,49,48,37,159,539,0,0,9,0,46,29,0,0,0,7,9,0,54,7,0,130,0,13,181,0,0,27
13,192.168.107.112,1693,73,194,4,1,115,691,125,44,0,7,0,0,0,80,324,26,44,0,177,359,0,0,0,0,90,46,0,0,0,0,0,0,35,11,0,108,0,3,99,2,0,40
74,192.168.107.169,1671,155,122,9,0,116,753,84,16,17,48,0,0,14,147,555,45,33,9,227,595,0,0,10,0,121,45,0,0,0,0,0,0,60,0,0,165,0,13,137,1,1,23
185,192.168.107.86,1659,113,73,0,0,78,737,71,54,2,28,6,1,0,95,334,39,51,4,284,511,0,1,33,10,87,15,1,0,0,0,0,0,40,0,0,158,0,3,185,3,0,8
120,192.168.107.210,1621,192,137,21,7,139,621,100,36,0,29,11,9,0,52,310,58,54,21,136,446,8,0,16,0,98,53,0,0,0,0,2,0,52,0,0,107,0,11,172,22,0,1
158,192.168.107.59,1601,105,147,6,30,51,562,122,43,11,8,9,0,3,20,406,28,7,4,167,520,0,0,5,0,62,22,17,0,0,0,0,12,18,0,0,151,0,18,149,10,0,47
163,192.168.107.64,1578,148,150,19,0,44,745,101,51,8,15,0,0,0,114,479,56,52,10,274,492,5,1,1,0,153,25,0,0,0,1,0,0,46,0,0,191,0,19,148,5,0,16
65,192.168.107.16,1577,106,142,13,9,77,698,127,15,0,48,0,0,6,84,290,40,31,0,207,431,0,0,2,1,38,69,0,0,0,0,0,0,45,0,0,140,0,1,122,36,0,24
115,192.168.107.206,1572,168,121,37,0,79,672,90,42,0,14,4,1,6,66,352,51,40,5,218,552,0,0,4,0,81,18,0,0,0,12,0,0,97,0,0,251,0,4,140,11,0,24
80,192.168.107.174,1567,110,97,20,0,87,555,112,18,0,21,10,0,15,99,290,25,10,4,224,574,0,3,7,0,107,22,0,0,0,0,0,0,21,0,0,140,0,14,161,15,0,15
109,192.168.107.200,1565,80,108,37,0,86,676,80,43,0,18,0,0,1,80,317,19,30,26,174,426,0,0,4,0,79,20,0,0,0,2,13,0,69,0,0,72,0,0,143,35,0,23
61,192.168.107.156,1565,111,202,4,9,100,726,129,72,0,14,0,0,0,118,314,67,63,0,268,666,1,0,1,0,68,25,0,0,0,0,0,0,38,0,0,139,0,38,124,14,0,42
56,192.168.107.151,1562,168,203,4,0,101,736,141,10,0,26,10,0,0,121,520,19,70,1,165,422,0,0,22,4,136,41,0,0,0,0,9,0,87,0,0,161,0,0,186,8,0,34
98,192.168.107.190,1551,122,217,23,0,136,726,99,35,4,27,1,5,4,89,362,97,49,15,243,523,0,0,6,0,77,86,0,0,0,0,0,0,52,0,0,119,0,19,147,20,0,24
135,192.168.107.36,1540,110,219,19,0,147,645,85,24,11,117,0,0,0,199,233,3,35,0,174,386,0,0,8,0,165,43,0,0,0,0,0,0,65,0,0,170,0,22,205,14,0,46
23,192.168.107.121,1535,96,92,5,2,82,668,55,16,0,46,0,18,0,81,243,24,38,1,153,448,4,0,1,0,78,36,0,0,0,0,0,0,58,1,0,185,0,11,206,0,0,5
153,192.168.107.54,1491,100,175,24,7,127,543,80,57,0,46,0,16,0,34,260,66,25,21,271,504,0,0,18,0,76,21,0,1,0,0,0,0,70,0,0,130,0,7,126,10,14,26
54,192.168.107.15,1486,109,144,12,1,87,692,90,78,0,80,7,0,2,75,423,57,40,18,265,439,13,0,4,0,85,74,2,0,0,0,0,0,53,0,0,188,0,9,127,12,0,33
133,192.168.107.34,1483,144,135,13,0,104,693,136,13,9,56,3,0,0,82,323,50,25,22,159,481,5,0,0,0,103,61,0,0,0,0,0,0,33,0,0,128,0,19,86,10,3,7
189,192.168.107.90,1455,72,182,21,0,117,790,112,32,0,42,20,0,0,112,355,58,35,15,180,414,0,0,3,0,43,48,0,0,0,0,0,0,60,0,0,213,0,4,143,30,0,32
11,192.168.107.110,1451,151,132,13,12,163,564,88,19,7,20,3,0,4,131,247,12,57,6,242,423,0,0,0,0,107,67,0,3,0,4,0,0,60,0,0,95,0,6,131,0,0,18
17,192.168.107.116,1435,110,142,7,0,66,522,68,35,0,17,16,8,0,141,314,31,37,13,156,515,0,0,42,0,83,48,0,0,0,0,0,0,74,0,0,128,0,4,172,8,2,9
182,192.168.107.83,1434,98,208,3,10,96,657,98,63,0,59,1,0,2,77,418,57,31,4,213,421,0,0,0,0,79,15,0,0,0,0,0,0,80,0,0,150,0,37,119,11,0,41
116,192.168.107.207,1431,127,102,56,4,78,626,84,43,0,39,1,0,2,84,343,5,26,8,194,423,0,5,11,0,46,10,0,0,0,0,11,0,39,0,0,137,0,0,87,19,0,9
60,192.168.107.155,1431,75,145,17,3,62,574,102,20,0,20,7,0,0,34,295,7,20,10,187,468,0,0,5,0,82,13,0,0,0,0,0,0,13,0,0,185,0,5,191,62,0,8
20,192.168.107.119,1393,117,130,0,4,84,525,41,47,0,15,6,0,2,74,278,26,5,3,178,350,0,0,1,0,70,3,0,2,0,0,0,0,33,0,0,126,0,4,161,7,0,6
82,192.168.107.176,1381,95,125,9,5,58,523,130,32,0,22,0,0,22,152,292,25,4,6,121,549,0,0,14,0,60,14,0,0,0,0,0,0,10,0,0,81,0,18,92,35,0,26
126,192.168.107.27,1381,161,69,2,0,118,623,91,23,4,40,2,6,0,98,308,45,33,6,190,407,0,0,1,0,62,21,0,0,0,0,0,0,81,0,0,181,0,7,113,6,0,28
66,192.168.107.160,1378,133,79,19,0,118,528,73,5,1,31,11,0,0,118,265,72,14,7,264,385,2,0,29,0,63,27,0,0,0,0,0,0,48,2,0,165,0,17,150,3,0,33
172,192.168.107.73,1371,79,89,32,7,108,522,77,14,8,13,0,0,2,22,223,47,15,14,179,462,0,0,8,0,84,49,0,0,0,0,0,0,75,0,0,186,0,0,109,30,0,17
165,192.168.107.66,1333,150,78,2,1,78,625,56,13,10,23,3,0,0,65,324,71,76,8,216,529,8,0,13,0,79,50,0,0,0,0,0,0,31,0,0,186,0,2,197,2,0,20
193,192.168.107.94,1318,94,127,9,4,119,405,104,11,0,17,5,0,0,111,297,51,28,2,169,374,0,3,27,0,88,29,0,0,0,0,0,0,9,0,0,92,0,1,153,10,0,14
15,192.168.107.114,1298,45,146,35,0,98,550,98,25,0,14,0,0,2,74,312,9,11,13,133,325,0,0,0,0,57,4,0,0,0,0,0,0,37,0,0,101,0,38,78,2,0,9
14,192.168.107.113,1280,37,115,16,0,50,501,60,13,9,29,0,0,0,97,375,11,27,5,164,509,0,0,18,0,59,26,0,0,0,0,0,0,46,6,0,151,0,3,85,7,0,14
142,192.168.107.43,1258,32,103,2,6,98,503,48,14,1,1,7,0,4,15,268,42,39,10,139,365,0,0,7,0,30,47,0,0,0,0,15,0,24,0,0,91,0,31,109,12,0,16
37,192.168.107.134,1256,38,153,10,0,71,530,85,5,0,43,0,2,0,27,253,12,62,0,112,320,0,0,1,0,63,42,0,0,0,0,0,0,57,0,0,100,0,10,138,0,0,57
67,192.168.107.161,1253,88,73,16,2,81,461,99,11,0,7,0,0,0,97,318,22,5,3,94,282,0,0,12,0,50,19,0,0,0,0,0,0,17,0,0,133,0,4,132,29,0,10
12,192.168.107.111,1253,49,81,5,2,69,398,86,27,0,6,3,0,0,33,283,29,45,14,120,241,1,0,0,0,67,24,0,0,0,0,0,0,40,1,0,73,0,11,63,2,0,12
170,192.168.107.71,1238,102,143,5,27,54,556,69,17,0,44,0,2,0,73,240,3,38,7,128,401,0,0,8,0,80,18,0,2,0,0,0,0,71,0,5,126,0,19,241,8,0,25
149,192.168.107.50,1210,125,64,20,0,62,556,124,7,0,40,2,0,0,45,341,52,38,11,194,363,0,0,4,0,70,31,0,0,0,0,4,0,52,0,0,80,0,0,123,18,0,7
38,192.168.107.135,1188,89,138,19,3,115,687,47,27,0,26,0,2,0,78,420,5,16,4,161,366,0,0,9,0,69,34,0,0,0,0,0,0,50,0,0,122,0,0,137,0,0,18
83,192.168.107.177,1184,50,40,22,0,22,441,50,7,0,8,3,21,0,38,273,25,17,9,168,300,0,0,5,0,15,44,0,0,3,0,0,0,26,0,0,58,0,5,160,7,0,1
188,192.168.107.89,1178,85,117,0,12,62,347,99,10,4,13,0,17,0,53,254,36,3,9,157,341,0,0,1,0,69,37,0,0,0,0,0,0,11,0,6,104,0,7,93,0,0,2
69,192.168.107.163,1170,86,103,12,0,83,581,72,16,4,50,0,0,0,49,221,28,29,7,239,343,10,0,0,0,67,18,0,0,0,0,0,0,52,0,0,133,0,10,109,3,0,2
132,192.168.107.33,1141,116,75,0,3,75,473,59,17,1,35,0,0,0,23,232,16,26,17,141,326,0,0,11,0,50,20,0,0,0,6,1,0,21,0,0,131,0,0,128,1,0,34
123,192.168.107.24,1130,85,63,0,0,40,326,131,17,0,8,4,0,0,37,216,49,24,16,74,282,7,0,7,0,76,47,0,0,0,2,0,0,43,0,0,89,0,43,135,2,0,8
27,192.168.107.125,1102,70,36,3,0,70,480,22,10,0,5,0,0,3,33,347,2,20,4,143,286,0,0,10,0,76,2,0,0,0,3,0,0,52,0,0,96,0,1,64,9,0,12
127,192.168.107.28,1094,109,61,20,0,100,635,114,13,0,10,0,1,0,56,263,19,23,25,195,304,0,0,0,0,54,6,16,0,0,0,0,18,18,0,0,116,0,0,122,6,0,10
76,192.168.107.170,1086,102,105,15,5,79,430,65,1,0,14,0,0,0,37,265,15,52,22,115,280,0,0,0,0,57,19,0,0,0,0,0,0,38,1,0,94,0,3,72,18,0,35
87,192.168.107.180,1069,104,105,2,3,63,488,108,19,0,26,10,0,0,49,211,32,22,0,200,433,7,0,3,0,53,4,0,0,0,0,2,0,49,5,0,114,0,0,105,14,0,18
176,192.168.107.77,1048,95,70,2,0,95,676,83,2,9,35,0,0,20,29,290,26,5,16,133,417,0,0,23,0,33,16,0,0,0,0,0,0,75,1,0,107,0,3,99,20,0,23
28,192.168.107.126,1043,94,77,0,1,36,530,57,32,0,37,3,0,0,67,280,8,26,12,151,480,0,0,1,0,65,15,0,0,0,0,0,0,50,0,0,197,0,8,120,12,0,27
84,192.168.107.178,1042,67,158,11,0,35,352,57,35,0,19,0,0,0,70,206,62,14,8,120,410,0,0,34,0,102,27,0,0,0,0,0,0,22,0,0,117,0,6,155,5,0,5
34,192.168.107.131,1033,75,107,15,0,43,428,46,27,8,25,0,0,0,60,299,20,33,0,72,289,0,0,12,0,46,14,0,0,0,0,0,0,39,0,0,132,0,3,83,12,0,35
63,192.168.107.158,1023,68,31,4,0,26,480,39,33,0,13,12,0,3,35,249,17,35,26,225,395,0,0,0,0,94,29,7,0,0,0,6,0,42,0,0,130,0,6,105,6,0,14
58,192.168.107.153,1009,108,73,12,1,59,377,57,20,0,13,16,1,2,77,277,26,7,7,114,280,0,0,20,0,23,18,0,0,0,0,0,0,20,0,0,68,0,19,147,8,0,5
48,192.168.107.144,1001,64,98,0,0,48,470,61,16,0,26,0,5,0,37,233,14,19,38,113,334,0,0,0,0,46,16,0,0,0,0,0,0,20,0,0,55,0,0,158,4,0,13
57,192.168.107.152,968,73,95,11,9,40,524,62,18,0,17,0,0,0,61,245,45,23,5,129,398,0,0,0,0,52,19,0,0,0,0,8,0,36,0,0,102,0,20,147,6,0,20
49,192.168.107.145,961,56,154,0,0,75,436,54,26,22,6,0,0,0,62,283,9,0,2,205,344,0,0,1,0,47,10,0,0,13,0,2,0,37,0,0,122,0,10,58,1,0,15
187,192.168.107.88,945,71,109,8,15,80,334,81,17,2,8,4,0,4,60,183,26,12,9,127,360,5,0,1,0,30,9,3,0,0,0,0,0,22,0,0,104,0,3,99,0,0,11
154,192.168.107.55,938,48,73,8,0,92,528,36,25,0,21,0,0,11,61,285,24,47,3,205,322,0,0,9,0,55,5,0,0,0,0,0,0,69,0,0,124,0,0,46,0,0,0
162,192.168.107.63,938,118,110,14,0,89,526,47,5,0,36,0,0,0,70,239,60,69,0,204,348,0,0,10,0,71,40,0,0,0,0,0,0,27,0,0,149,0,1,96,5,0,16
16,192.168.107.115,877,85,64,1,0,57,375,43,13,0,5,2,0,0,58,204,29,29,46,125,322,0,0,4,0,86,22,0,0,0,0,0,0,32,0,0,102,0,2,118,13,0,11
5,192.168.107.105,861,50,66,10,0,59,469,109,4,0,21,0,0,0,32,184,57,12,3,82,238,0,0,7,0,24,16,0,0,0,0,0,0,75,0,0,102,0,0,123,1,0,2
97,192.168.107.19,847,58,120,15,0,53,319,27,29,0,41,0,0,0,50,148,22,15,3,117,205,0,0,19,0,50,27,0,0,0,0,0,0,20,0,0,99,0,0,101,14,0,11
94,192.168.107.187,832,118,51,39,1,61,265,24,27,0,22,0,0,0,77,147,4,2,5,58,198,0,0,0,0,51,10,0,0,0,0,0,0,30,3,0,79,0,3,54,11,0,6
31,192.168.107.129,802,32,82,3,11,31,352,53,32,0,2,0,0,0,32,193,17,38,7,107,267,3,0,19,0,40,21,0,0,0,0,0,0,35,0,0,84,0,18,57,8,0,0
0,192.168.107.100,778,94,51,4,0,33,294,94,9,0,17,0,0,1,60,215,42,13,8,113,317,0,0,0,0,35,30,0,0,0,0,0,0,34,0,0,65,0,0,85,1,0,40
186,192.168.107.87,747,36,82,0,0,119,390,35,32,0,8,0,0,0,29,191,22,4,5,131,195,0,0,3,0,36,28,0,0,0,0,0,0,10,0,0,97,9,9,104,0,0,34
52,192.168.107.148,723,41,60,14,7,57,218,28,10,0,10,8,0,0,52,127,6,21,2,88,184,0,0,1,0,12,35,0,0,0,0,0,0,10,0,0,73,0,4,73,7,0,20
181,192.168.107.82,718,88,62,21,1,57,313,77,8,0,20,0,0,11,28,121,12,6,4,86,161,0,0,0,0,79,21,0,0,0,0,0,0,19,0,0,48,0,6,109,0,0,4
110,192.168.107.201,709,37,74,8,0,62,296,43,8,0,14,0,0,9,67,128,39,25,8,102,223,0,0,2,0,29,24,0,0,0,0,0,0,78,0,0,35,0,3,77,18,0,11
122,192.168.107.23,684,25,90,7,0,55,290,3,1,17,10,3,1,0,11,161,10,28,1,65,170,0,0,0,0,16,17,0,0,0,0,0,0,37,0,0,90,0,25,43,7,0,25
90,192.168.107.183,670,47,66,0,0,39,455,82,13,0,28,0,0,0,29,197,23,3,1,105,270,0,0,4,0,48,43,0,0,0,0,0,0,10,0,0,71,0,3,73,1,0,6
99,192.168.107.191,565,26,30,0,0,112,235,46,2,0,26,0,0,0,23,184,3,2,6,21,170,0,0,23,0,48,17,0,0,0,0,0,0,7,0,0,40,0,2,71,0,0,2
79,192.168.107.173,561,26,63,0,0,24,311,8,19,5,51,12,0,3,29,173,21,6,2,63,123,0,0,0,0,22,9,0,0,0,0,0,0,31,0,0,83,0,0,19,0,0,7
25,192.168.107.123,523,35,42,0,5,36,236,42,1,4,10,0,0,11,20,149,4,12,0,60,176,0,0,0,0,56,15,0,0,0,1,0,0,10,0,0,29,0,0,79,4,0,8
108,192.168.107.20,521,20,23,20,0,28,186,24,11,0,3,0,0,0,59,89,19,16,0,21,148,0,0,14,0,19,10,0,0,0,0,0,0,27,0,0,43,0,0,60,3,0,16
166,192.168.107.67,517,33,91,9,0,41,210,24,7,1,7,0,7,0,67,196,4,8,0,79,364,0,0,9,0,70,23,0,0,0,0,0,0,8,0,0,94,0,9,67,0,0,4
2,192.168.107.102,510,17,31,0,0,59,159,28,0,8,10,4,0,0,1,128,15,0,0,93,141,0,0,1,0,23,19,0,0,0,0,0,0,53,0,0,26,0,1,41,1,0,3
6,192.168.107.106,506,30,32,3,0,56,213,39,0,0,18,0,0,0,10,111,8,13,11,100,170,0,0,0,0,29,9,0,0,0,0,0,0,25,0,0,73,0,12,38,8,0,1
86,192.168.107.18,495,14,14,0,1,43,164,36,3,8,0,11,0,0,14,94,25,1,7,118,139,0,0,0,0,18,3,0,0,0,0,0,0,44,0,0,22,0,18,35,14,0,8
156,192.168.107.57,437,25,30,0,0,53,127,7,27,0,12,0,0,8,13,136,9,10,0,38,141,0,0,3,0,45,12,0,0,0,0,0,0,8,0,0,44,0,16,62,4,0,0
51,192.168.107.147,410,13,7,3,0,30,271,25,1,0,1,10,0,0,12,115,18,0,0,31,136,0,0,10,0,10,2,0,0,0,0,0,0,31,0,0,57,0,4,5,6,0,1
24,192.168.107.122,401,36,59,0,0,20,156,62,10,0,0,0,0,0,2,82,13,27,0,33,105,3,0,0,0,3,8,0,0,0,0,0,0,24,0,0,49,0,0,8,0,0,0
46,192.168.107.142,398,15,54,8,0,5,140,7,6,0,25,0,4,0,12,82,2,4,2,36,99,0,0,0,0,19,7,0,0,0,0,0,0,10,0,0,18,0,0,53,0,0,8
113,192.168.107.204,373,16,54,0,10,22,108,5,17,0,6,0,0,0,21,75,0,6,0,68,101,0,0,6,0,22,17,0,0,11,3,0,0,26,0,0,22,0,0,3,1,0,4
73,192.168.107.168,367,4,18,0,0,21,165,51,16,0,10,0,0,0,16,81,0,25,0,44,114,0,0,0,0,43,2,0,0,0,0,0,0,41,0,0,34,0,2,12,17,0,9
8,192.168.107.108,357,16,9,0,24,13,114,17,6,0,9,0,0,0,14,63,24,0,0,48,69,0,0,0,0,9,4,0,0,0,0,1,0,0,0,0,41,0,0,54,0,0,0
45,192.168.107.141,353,34,50,0,0,10,224,34,30,0,16,0,0,0,44,50,0,6,0,77,153,0,0,7,0,10,22,0,0,0,0,0,0,13,0,0,63,0,9,47,12,0,11
68,192.168.107.162,344,16,35,0,0,30,152,9,7,0,3,0,0,0,21,77,10,2,0,40,161,0,0,0,0,23,3,0,0,0,0,0,0,9,0,0,58,0,0,21,0,0,0
198,192.168.107.99,276,37,53,0,12,24,139,10,6,2,8,0,0,0,7,76,3,5,0,53,147,0,0,0,0,14,11,0,0,0,0,0,0,23,0,0,9,0,4,20,0,0,1
121,192.168.107.22,236,31,1,0,0,11,78,8,0,8,0,0,0,0,0,27,0,15,2,5,42,0,0,0,0,2,17,0,0,0,0,0,0,0,0,0,0,0,0,10,0,0,6
180,192.168.107.81,225,17,23,2,0,17,87,15,0,0,0,0,0,0,8,30,0,0,10,16,87,0,0,0,0,27,0,0,0,0,0,0,0,1,0,0,17,0,0,7,1,0,7
196,192.168.107.97,203,7,7,0,0,3,82,4,3,0,0,6,0,0,4,39,0,3,0,42,105,0,0,3,0,8,12,0,0,0,0,0,0,0,0,0,16,0,0,15,0,0,8
47,192.168.107.143,67,4,3,0,0,11,40,0,3,0,0,0,0,0,0,12,0,0,9,3,18,0,0,0,0,0,4,0,0,0,0,0,0,6,0,0,0,0,0,28,0,0,0
